`define KIWI